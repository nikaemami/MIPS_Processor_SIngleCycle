module datapath(MD_out, sel_wr_2, sel_wr_1, RegWrite, sel_B, ALU_control, MemtoReg, branch, sel_data, sel_pc_1, pc_src, clk, rst, inst_out, slt_sel, alu_out, pc_out, Read2);
	input [31:0] inst_out, MD_out;
	input [2:0] ALU_control;
	input sel_wr_2, sel_wr_1, RegWrite, sel_B, MemtoReg, branch, sel_data, sel_pc_1, pc_src, clk, rst, slt_sel;
	output [31:0] alu_out, pc_out, Read2;
	wire [31:0] inst_out, shl_out, M1_out, Read1, Read2, add1_out, MemtoReg_out, SE_out, M2_out;
	wire [31:0] M9_out ,M10_out ,M5_out ,M4_out ,adder2_out ,shl2_out ,MD_out, alu_out, pc_src_out, pc_out; 
	wire [4:0] M7_out, M8_out;
	wire zero, sel_M4, negative;
	assign sel_M4 = zero & branch;
	Sign_Extend SE(inst_out[15:0], SE_out);
	Sign_extend_26 SE26(inst_out[25:0], shl_out);
	Shift_Left_2 SHL2(SE_out, shl2_out);
	adder_32 adder1(pc_out, {32'd4}, add1_out);
	adder_32 adder2(add1_out, shl2_out, adder2_out);
	Register_File RF(clk, rst, inst_out[25:21], inst_out[20:16], M8_out, M10_out, RegWrite, Read1, Read2);
	ALU alu(Read1, M2_out, ALU_control, alu_out, zero, negative);
	PC pc(clk, rst, pc_src_out, pc_out);
	mux2to1_32 M1(add1_out, MemtoReg_out, sel_data, M1_out);
	mux2to1_32 M2(Read2, SE_out, sel_B, M2_out);
	mux2to1_32 M3(alu_out, MD_out, MemtoReg, MemtoReg_out);
	mux2to1_32 M4(add1_out, adder2_out, sel_M4, M4_out);
	mux2to1_32 M5(Read1, shl_out, sel_pc_1, M5_out);
	mux2to1_32 M6(M4_out, M5_out, pc_src, pc_src_out);
	mux2to1_32 M9({32'd0}, {32'd1}, negative, M9_out);
	mux2to1_32 M10(M1_out, M9_out, slt_sel, M10_out);
	mux2to1_5 M7(inst_out[20:16], inst_out[15:11], sel_wr_2, M7_out);
	mux2to1_5 M8(M7_out, {5'd31}, sel_wr_1, M8_out);
endmodule
